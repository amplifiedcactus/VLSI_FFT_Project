//FFT Module

//State machine:
//Idle State
//Retrieve data from RAM State, put it in the cache
//Computing FFT stage 1
//Computing FFT stage 2
//Computing FFT stage 3
//Computing FFT stage 4
//Send results to RAM State

//Define twiddle factor registers

//Define registers for storing results of each stage (cache)

//For each stage, instantiate a FFTStage module with the correct inputs (from storage registers), and connect the outputs to the cache


