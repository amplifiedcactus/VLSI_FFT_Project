//Module that takes 8 pairs of 32 bit complex numbers (16 total) and uses the MultiplyAddUnit module to compute a single stage of a 16-point FFT 
module FFTStage(inputVector, outputVector, Clk, Rst)

endmodule