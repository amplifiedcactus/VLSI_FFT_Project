//Module that takes 3 32 bit complex numbers as inputs, A, B and w. 2 32 bit complex numbers are output, Y and Z.
//Y is set equal to A+(B*w)
//Z is set equal to A-(B*w)
module MultiplyAddUnit (A, B, w, Y, Z, Clk, Rst)

endmodule